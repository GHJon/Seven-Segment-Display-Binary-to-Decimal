LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

Entity RODR_MASTERMAP IS
	PORT(RODR_SIGBIT      : IN STD_LOGIC;
			  RODR_IN       : IN STD_LOGIC_VECTOR (7 downto 0) ;
			  RODR_ONES     : OUT STD_LOGIC_VECTOR (6 downto 0);
			  RODR_TENS     : OUT STD_LOGIC_VECTOR (6 downto 0);
			  RODR_HUNDREDS : OUT STD_LOGIC_VECTOR (6 downto 0);
			  RODR_SIGN		 : OUT STD_LOGIC_VECTOR (6 downto 0);
			  RODR_LEDONOFF : OUT STD_LOGIC_VECTOR (8 downto 0);
			  RODR_DISP4     : OUT STD_LOGIC_VECTOR (6 downto 0);
			  RODR_DISP5     : OUT STD_LOGIC_VECTOR (6 downto 0);
			  RODR_DISP6     : OUT STD_LOGIC_VECTOR (6 downto 0);
			  RODR_DISP7     : OUT STD_LOGIC_VECTOR (6 downto 0));


END RODR_MASTERMAP;

ARCHITECTURE CONNECTIONS of RODR_MASTERMAP IS
	Component RODR_UnsignedSigned IS
		PORT(RODR_SIGBIT : IN STD_LOGIC;
			RODR_IN   : IN STD_LOGIC_VECTOR (7 downto 0) ;
			RODR_OUT  : OUT STD_LOGIC_VECTOR (7 downto 0);
			RODR_LEDS : OUT STD_LOGIC_VECTOR (8 downto 0));		
	END Component;

	Component RODR_BINARYBCD
		PORT(RODR_IN: IN STD_LOGIC_VECTOR (7 downto 0) ;
		   RODR_OUT : OUT STD_LOGIC_VECTOR (11 downto 0));
	END Component ;

	Component RODR_BCDDecoder
		PORT(RODR_IN: IN STD_LOGIC_VECTOR (3 downto 0) ;
	      RODR_OUT : OUT STD_LOGIC_VECTOR (6 downto 0));
	END Component ;
	
	Component RODR_PlusMinus
	PORT(RODR_SIGBIT : IN STD_LOGIC;
		  RODR_IN: IN STD_LOGIC_VECTOR (7 downto 0);
	     RODR_OUT : OUT STD_LOGIC_VECTOR (6 downto 0));
	END Component;
	
	Component RODR_NOOUTPUT
			PORT(RODR_OUT : OUT STD_LOGIC_VECTOR (6 downto 0));
	END Component ;
	
signal RODR_TCO : STD_LOGIC_VECTOR (7 downto 0);		--TCO = TWo's Complement Output
signal RODR_BCD : STD_LOGIC_VECTOR (11 downto 0);
signal RODR_BCD_ONE : STD_LOGIC_VECTOR (3 downto 0);
signal RODR_BCD_TEN : STD_LOGIC_VECTOR (3 downto 0);
signal RODR_BCD_HUNDRED : STD_LOGIC_VECTOR (3 downto 0);

BEGIN
	
	RODR_TWOSCOMPLEMENT   : RODR_UnsignedSigned  PORT MAP(RODR_SIGBIT, RODR_IN, RODR_TCO, RODR_LEDONOFF);
	RODR_BINARYTOBCD      : RODR_BINARYBCD 		PORT MAP(RODR_TCO, RODR_BCD);
	
	RODR_BCD_ONE <= STD_LOGIC_VECTOR (RODR_BCD(3 downto 0));
	RODR_BCD_TEN <= STD_LOGIC_VECTOR (RODR_BCD(7 downto 4));
	RODR_BCD_HUNDRED <= STD_LOGIC_VECTOR (RODR_BCD(11 downto 8));
	
	
	RODR_DecoderONES 		 : RODR_BCDDecoder 		PORT MAP(RODR_BCD_ONE, RODR_ONES);
	RODR_DecoderTENS		 : RODR_BCDDecoder 		PORT MAP(RODR_BCD_TEN, RODR_TENS);
	RODR_DecoderHUNDREDS  : RODR_BCDDecoder 		PORT MAP(RODR_BCD_HUNDRED, RODR_HUNDREDS);
	RODR_POSNEG				 : RODR_PlusMinus			PORT MAP (RODR_SIGBIT, RODR_IN, RODR_SIGN);
	RODR_DISPLAYOFF4			 : RODR_NOOUTPUT			PORT MAP (RODR_DISP4);
	RODR_DISPLAYOFF5			 : RODR_NOOUTPUT			PORT MAP (RODR_DISP5);
	RODR_DISPLAYOFF6			 : RODR_NOOUTPUT			PORT MAP (RODR_DISP6);
	RODR_DISPLAYOFF7			 : RODR_NOOUTPUT			PORT MAP (RODR_DISP7);

END CONNECTIONS;